////////////////////////////////////////////////////////////////////////////////
//                                                                            //
// Copyright 2025 ETH Zurich and University of Bologna.                       //
// Copyright and related rights are licensed under the Solderpad Hardware     //
// License, Version 0.51 (the "License"); you may not use this file except in //
// compliance with the License.  You may obtain a copy of the License at      //
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law  //
// or agreed to in writing, software, hardware and materials distributed under//
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR     //
// CONDITIONS OF ANY KIND, either express or implied. See the License for the //
// specific language governing permissions and limitations under the License. //
//                                                                            //
//                                                                            //
// Engineer:      Maurus Item - itemm@student.ethz.ch                         //
//                                                                            //
// Additional contributions by:                                               //
//                                                                            //
//                                                                            //
//                                                                            //
// Create Date:    02/01/2025                                                 //
// Design Name:    redundant shared fpu cluster                               //
// Module Name:    fpu_demux                                                  //
// Project Name:   Redundant Floating-Point Units and Accelerators            //
// Language:       SystemVerilog                                              //
//                                                                            //
// Description:                                                               //
// This module demuxes the FPU and the shared Division without any statefull  //
// behaviour and is as such stall-safe. Cores using it need to deal with      //
// out-of-order results themselves!                                           //
//                                                                            //
// Revision:                                                                  //
// Revision v0.1 - 02/01/2025 : File Created                                  //
//                                                                            //
// Additional Comments:                                                       //
//                                                                            //
//                                                                            //
//                                                                            //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////

module fpu_demux
#(
    parameter DATA_WIDTH         = 32,
    parameter FP_TYPE_WIDTH      = 5,
    parameter NB_CORE_ARGS       = 3,
    parameter CORE_OPCODE_WIDTH  = 6,
    parameter CORE_DSFLAGS_CPU   = 15,
    parameter CORE_USFLAGS_CPU   = 5,

    parameter NB_APU_ARGS        = 3,
    parameter APU_OPCODE_WIDTH   = 6,
    parameter APU_DSFLAGS_CPU    = 15,
    parameter APU_USFLAGS_CPU    = 5,

    parameter NB_FPNEW_ARGS      = 3,
    parameter FPNEW_OPCODE_WIDTH = 6,
    parameter FPNEW_DSFLAGS_CPU  = 15,
    parameter FPNEW_USFLAGS_CPU  = 5,

    parameter APU_ID             = 1,
    parameter FPNEW_ID           = 0
)
(
    input  logic                                         clk,
    input  logic                                         rst_n,

    // CORE SIDE: Slave port
    // request channel
    input  logic                                         core_slave_req_i,
    output logic                                         core_slave_gnt_o,
    input  logic [FP_TYPE_WIDTH-1:0]                     core_slave_type_i,
    input  logic [NB_CORE_ARGS-1:0][DATA_WIDTH-1:0]      core_slave_operands_i,
    input  logic [CORE_OPCODE_WIDTH-1:0]                 core_slave_op_i,
    input  logic [CORE_DSFLAGS_CPU-1:0]                  core_slave_flags_i,
    // response channel
    input  logic                                         core_slave_rready_i,
    output logic                                         core_slave_rvalid_o,
    output logic [DATA_WIDTH-1:0]                        core_slave_rdata_o,
    output logic [CORE_USFLAGS_CPU-1:0]                  core_slave_rflags_o,

    // APU Side: Master port
    // request channel
    output logic                                         apu_req_o,
    input  logic                                         apu_gnt_i,
    output logic [NB_APU_ARGS-1:0][DATA_WIDTH-1:0]       apu_operands_o,
    output logic [APU_OPCODE_WIDTH-1:0]                  apu_op_o,
    output logic [APU_DSFLAGS_CPU-1:0]                   apu_flags_o,
    // response channel
    output logic                                         apu_rready_o,
    input  logic                                         apu_rvalid_i,
    input  logic [DATA_WIDTH-1:0]                        apu_rdata_i,
    input  logic [APU_USFLAGS_CPU-1:0]                   apu_rflags_i,

    // FPNEW Side: Master port
    // request channel
    output logic                                         fpnew_req_o,
    input  logic                                         fpnew_gnt_i,
    output logic [NB_FPNEW_ARGS-1:0][DATA_WIDTH-1:0]     fpnew_operands_o,
    output logic [FPNEW_OPCODE_WIDTH-1:0]                fpnew_op_o,
    output logic [FPNEW_DSFLAGS_CPU-1:0]                 fpnew_flags_o,
    // response channel
    output logic                                         fpnew_rready_o,
    input  logic                                         fpnew_rvalid_i,
    input  logic [DATA_WIDTH-1:0]                        fpnew_rdata_i,
    input  logic [FPNEW_USFLAGS_CPU-1:0]                 fpnew_rflags_i
);  
    
    // Non-handshake stuff gets wired straight through
    assign fpnew_operands_o = core_slave_operands_i[NB_FPNEW_ARGS-1:0];
    assign fpnew_op_o       = core_slave_op_i[FPNEW_OPCODE_WIDTH-1:0];
    assign fpnew_flags_o    = core_slave_flags_i[FPNEW_DSFLAGS_CPU-1:0];

    assign apu_operands_o   = core_slave_operands_i[NB_APU_ARGS-1:0];
    assign apu_op_o         = core_slave_op_i[APU_OPCODE_WIDTH-1:0];
    assign apu_flags_o      = core_slave_flags_i[APU_DSFLAGS_CPU-1:0];

    // Input Handshake according to select signal
    always_comb begin
        apu_req_o        = 1'b0;
        fpnew_req_o      = 1'b0;     
        core_slave_gnt_o = 1'b0;    

        case (core_slave_type_i)
            APU_ID: begin
                apu_req_o         = core_slave_req_i;
                core_slave_gnt_o  = apu_gnt_i;
            end

            FPNEW_ID: begin
                fpnew_req_o       = core_slave_req_i;
                core_slave_gnt_o  = fpnew_gnt_i;
            end

            /* add other mux outputs here in the same format */
        endcase
    end

    // Output Handshake according to valid, prioritizing fpu inputs
    always_comb begin
        core_slave_rvalid_o   = fpnew_rvalid_i | apu_rvalid_i;
        fpnew_rready_o = 1'b0;
        apu_rready_o = 1'b0;

        if (fpnew_rvalid_i) begin
            fpnew_rready_o       = core_slave_rready_i;
            core_slave_rdata_o   = fpnew_rdata_i;
            core_slave_rflags_o  = fpnew_rflags_i; 

        /* add other mux inputs here in the same format with else if */
 
        end else begin
            apu_rready_o         = core_slave_rready_i;
            core_slave_rdata_o   = apu_rdata_i;
            core_slave_rflags_o  = apu_rflags_i;
        end
    end

endmodule